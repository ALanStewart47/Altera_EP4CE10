module top_led(
    input       sys_clk,
    input       sys_rst_n,

    input       key,
    output      led
);

wire key_value;
wire key_flag;


key_fliter  u_key_fliter(
    
);